module instmemory( write, addr, datain, dataout, clk, reset);
	input [31:0] datain;
	input [15:0] addr;
	input write, clk, reset;
	output [31:0] dataout;
	
	reg[31:0] mem[255 : 0];
	
	assign dataout = mem[addr];
	
	always @(posedge clk) begin
		if(reset) begin
			mem[0] <=32'b0110111101111010_0000000000001010;
			mem[1] <=32'b1101100000111011_1100000000000000;
			mem[2] <=32'b0110111100111000_0000000000000010;
			mem[3] <=32'b1000111101000000_0000000000000010;
			mem[4] <=32'b0110111101111011_1111111111111110;
			mem[5] <=32'b0110100000000000_0000000000000000;
			mem[6] <=32'b0110111110111100_0000000000001010;
			mem[7] <=32'b0110100001000010_0000000000001010;
			mem[8] <=32'b0101000010000000_0000000000000000;
			mem[9] <=32'b0110100010000100_0000000000000110;
			mem[10] <=32'b0101000011000000_0000000000000000;
			mem[11] <=32'b0110100011000110_0000000000001000;
			mem[12] <=32'b0101100100000101_1110000000000000;
			mem[13] <=32'b0101100101000111_1110000000000000;
			mem[14] <=32'b0100000110001010_0100000000000000;
			mem[15] <=32'b1000000000001100_0000000000100110;
			mem[16] <=32'b0000100000000000_0000000000000000;
			mem[17] <=32'b1101100000000110_0100000000000000;
			mem[18] <=32'b1101100000000100_0101000000000000;
			mem[19] <=32'b0110100011000111_1111111111111110;
			mem[20] <=32'b0110100010000101_1111111111111110;
			mem[21] <=32'b1000100011000000_0000000000011000;
			mem[22] <=32'b0000100000000000_0000000000000000;
			mem[23] <=32'b0110100001000011_1111111111111110;
			mem[24] <=32'b1000100000000010_0000000000010000;
			mem[25] <=32'b0101011101000000_0000000000000000;
			mem[26] <=32'b0101011100000000_0000000000000000;
			mem[27] <=32'b0110111101111010_0000000000001010;
			mem[28] <=32'b0101100100111001_1110000000000000;
			mem[29] <=32'b0110111101111011_1111111111111110;
			mem[30] <=32'b0110111100111000_0000000000000010;
			mem[31] <=32'b1000111101000000_0000000000111000;
		end
		else begin
			if(write==1)
				mem[addr]<=datain;
			
		end

	end
endmodule
