module datamemory( write, addr, datain, dataout, clk, reset);
	input [31:0] datain;
	input [15:0] addr;
	input write, clk, reset;
	output reg[31:0] dataout;
	
	reg[31:0] mem[255 : 0];
	
	always @(posedge clk) begin
		if(reset) begin
			mem[0] <=32'b0000000000000000_0000000000000000;
			mem[1] <=32'b0000000000000000_0000000000000000;
			mem[2] <=32'b0000000000000000_0000000000000000;
			mem[3] <=32'b0000000000000000_0000000000000000;
			mem[4] <=32'b0000000000000000_0000000000000000;
			mem[5] <=32'b0000000000000000_0000000000000000;
			mem[6] <=32'b0000000000000000_0000000000000000;
			mem[7] <=32'b0000000000000000_0000000000000000;
			mem[8] <=32'b0000000000000000_0000000000000000;
			mem[9] <=32'b0000000000000000_0000000000000000;
			mem[10]<=32'b0000000000000000_0000000000000000;
			mem[11]<=32'b0000000000000000_0000000000000000;
			mem[12]<=32'b0000000000000000_0000000000000000;
			mem[13]<=32'b0000000000000000_0000000000000000;
			mem[14]<=32'b0000000000000000_0000000000000000;
			mem[15]<=32'b0000000000000000_0000000000000000;
			mem[16]<=32'b0000000000000000_0000000000000000;
			mem[17]<=32'b0000000000000000_0000000000000000;
			mem[18]<=32'b0000000000000000_0000000000000000;
			mem[19]<=32'b0000000000000000_0000000000000000;
			mem[20]<=32'b0000000000000000_0000000000000000;
			mem[21]<=32'b0000000000000000_0000000000000000;
			mem[22]<=32'b0000000000000000_0000000000000000;
			mem[23]<=32'b0000000000000000_0000000000000000;
			mem[24]<=32'b0000000000000000_0000000000000000;
			mem[25]<=32'b0000000000000000_0000000000000000;
			mem[26]<=32'b0000000000000000_0000000000000000;
			mem[27]<=32'b0000000000000000_0000000000000000;
			mem[28]<=32'b0000000000000000_0000000000000000;
			mem[29]<=32'b0000000000000000_0000000000000000;
			mem[30]<=32'b0000000000000000_0000000000000000;
			mem[31]<=32'b0000000000000000_0000000000000000;
			mem[32]<=32'b0000000000000000_0000000000000000;
		end
		else begin
			if(write==1)
				mem[addr]<=datain;
			dataout<= mem[addr];
		end

	end
endmodule
