module instmemory( write, addr, datain, dataout, clk, reset);
	input [31:0] datain;
	input [15:0] addr;
	input write, clk, reset;
	output [31:0] dataout;
	
	reg[31:0] mem[255 : 0];
	
	assign dataout = mem[addr];
	
	always @(posedge clk) begin
		if(reset) begin
			mem[0] <=32'b0110111111111110_0000000000110110;
			mem[1] <=32'b0110100000000000_0000000000000000;
			mem[2] <=32'b0101000001000000_0000000000000000;
			mem[3] <=32'b0110100011000110_0000000000000110;
			mem[4] <=32'b0101000010000000_0000000000000000;
			mem[5] <=32'b0110100001000010_0000000000000110;
			mem[6] <=32'b0110100010000100_0000000000000110;
			mem[7] <=32'b0110100001000011_1111111111111110;
			mem[8] <=32'b0110100010000101_1111111111111110;
			mem[9] <=32'b0100111110001000_0011000010000000;
			mem[10] <=32'b0101000101000000_0000000000000000;
			mem[11] <=32'b0000100101001010_0010000000000000;
			mem[12] <=32'b0101001101000000_0000000000000000;
			mem[13] <=32'b0000101101011010_0100000000000000;
			mem[14] <=32'b0000101101011010_0101000000000000;
			mem[15] <=32'b0110101101011010_0000000000100100;
			mem[16] <=32'b0110100101001010_0000000000010010;
			mem[17] <=32'b0101000110000000_0000000000000000;
			mem[18] <=32'b0110100110001100_0000000000000100;
			mem[19] <=32'b0101000111000000_0000000000000000;
			mem[20] <=32'b0101101000111110_0100000000000000;
			mem[21] <=32'b0101101001111110_0101000000000000;
			mem[22] <=32'b0100111110011000_1000010010000000;
			mem[23] <=32'b0000100111001110_1100000000000000;
			mem[24] <=32'b0110100100001000_0000000000000010;
			mem[25] <=32'b0110100101001010_0000000000000110;
			mem[26] <=32'b1000100110000000_0000000000101000;
			mem[27] <=32'b0110100110001101_1111111111111110;
			mem[28] <=32'b1101100000011010_0111000000000000;
			mem[29] <=32'b1000100010000000_0000000000010000;
			mem[30] <=32'b0000100000000000_0000000000000000;
			mem[31] <=32'b1000100001000000_0000000000001100;
			mem[32] <=32'b0000100000000000_0000000000000000;
		end
		else begin
			if(write==1)
				mem[addr]<=datain;
			
		end

	end
endmodule
